
module max10clk (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
